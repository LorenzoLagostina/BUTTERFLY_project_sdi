library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
package bf is
	type stage is array (0 to 15) of signed(19 downto 0);
end bf;
